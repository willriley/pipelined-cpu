module pipelined_cpu(input CLOCK_50);



endmodule